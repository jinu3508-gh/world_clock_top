`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/11/24 13:27:25
// Design Name: 
// Module Name: clock
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module world_clock_top(
    input clk,
    input rst,

    // ���� ��ư (1~7)
    input adj_min_btn,      // BTN 2 (�ð�: �� ���� / �˶�: �� ����)
    input adj_hour_btn,     // BTN 1 (�ð�: �� ���� / �˶�: �� ����)
    input mode_toggle_btn,  // BTN 3 (12/24H ���)
    input paris_btn,        // BTN 5 (������ 5�� -> Paris / Alarm 2)
    input ny_btn,           // BTN 4 (������ 4�� -> NY / Alarm 1)
    input uk_btn,           // BTN 6 (UK / Alarm 3)
    input korea_btn,        // BTN 7 (Korea)

    // �߰��� ��ư (8~10) - Ÿ�̸ӿ� (*, 0, #)
    input btn_tm_min,       // Key * (Ÿ�̸� �� / �˶� ����)
    input btn_tm_sec,       // Key 0 (Ÿ�̸� �� / �˶� ����)
    input btn_tm_start,     // Key # (Ÿ�̸� ���� / �˶� ����)
    
    // �˶� ���¿� ��ư (Key 8)
    input btn_num_8,

    // ����ġ
    input sw_timer,         // SW3 (Timer Mode)
    input sw_alarm,         // SW4 (Alarm Set Mode)

    // ���
    output [7:0] seg_data,
    output [7:0] seg_com,
    output LCD_E,
    output LCD_RS,
    output LCD_RW,
    output [7:0] LCD_DATA,
    output reg piezo,       // �ǿ��� ���
    
    // LED ���
    output wire tm_led_r, tm_led_g, tm_led_b, // Ÿ�̸� 3�� LED
    output wire alm_led1, alm_led2, alm_led3  // �˶� 1/2/3 ���� LED
);

    // ==================================================
    // 1. ��ư �Է� ó�� (Oneshot) - �� 11��
    // ==================================================
    wire [10:0] btn_trig; 

    // oneshot ����� �Է� ��Ʈ ������ �߿��մϴ�.
    oneshot_universal #(.WIDTH(11)) U_OS (
        .clk     (clk),
        .rst     (rst),
        .btn     ({btn_num_8, btn_tm_start, btn_tm_sec, btn_tm_min,
                    adj_min_btn, adj_hour_btn, mode_toggle_btn,
                    paris_btn,    ny_btn,       uk_btn, korea_btn}),
        .btn_trig(btn_trig)
    );

    // --- ��ư ��ȣ ���� (������ ��ư ����) ---
    
    // [Keypad]
    // [���� 1] Key 8��(btn_trig[10])�� ��ɺ��� �и�
    wire btn_key8_raw = btn_trig[10];

    // SW3(Timer)�� ���� ������ 'Ÿ�̸� ����', ���� ������ '�˶� ����'
    wire btn_timer_reset_p = (sw_timer) ? btn_key8_raw : 1'b0;
    wire btn_alarm_reset_p = (sw_timer) ? 1'b0 : btn_key8_raw;
    
    wire tm_start_p = btn_trig[9]; // Key #
    wire tm_sec_p   = btn_trig[8]; // Key 0
    wire tm_min_p   = btn_trig[7]; // Key *
    
    // �˶� �ð�(Alarm Clock)�� �︱ �� ���� ��ȣ (�� �� �ƹ��ų�)
    wire alarm_stop_signal = tm_start_p | tm_sec_p | tm_min_p;

    // [Time Control]
    wire adj_min_raw_p  = btn_trig[6]; // BTN 2
    wire adj_hour_raw_p = btn_trig[5]; // BTN 1
    wire mode_toggle_p  = btn_trig[4]; // BTN 3
    
    // [City Control]
    // oneshot �Է� ����: {..., paris_btn, ny_btn, ...}
    // btn_trig[3] = paris_btn (������ 5��)
    // btn_trig[2] = ny_btn    (������ 4��)
    
    wire btn_paris_raw = btn_trig[3]; // BTN 5
    wire btn_ny_raw    = btn_trig[2]; // BTN 4
    wire btn_uk_raw    = btn_trig[1]; // BTN 6
    wire btn_korea_raw = btn_trig[0]; // BTN 7

    
    // ==================================================
    // [��ư MUX ����] SW4 ���¿� ���� ��� �й�
    // ==================================================

    // 1. �ð� ���� (BTN 1, 2)
    // SW4 ON -> �˶� �ð� ����, SW4 OFF -> ���� �ð� ����
    wire time_adj_min_p   = (sw_alarm) ? 1'b0 : adj_min_raw_p;
    wire time_adj_hour_p  = (sw_alarm) ? 1'b0 : adj_hour_raw_p;
    
    wire alarm_adj_min_p  = (sw_alarm) ? adj_min_raw_p : 1'b0;
    wire alarm_adj_hour_p = (sw_alarm) ? adj_hour_raw_p : 1'b0;

    // 2. ���� ���� vs �˶� ���� ���� (BTN 4, 5, 6)
    
    // �ð� ���� (SW4 OFF): ���� ����
    wire clk_ny_p    = (sw_alarm) ? 1'b0 : btn_ny_raw;    // BTN 4 -> NY
    wire clk_paris_p = (sw_alarm) ? 1'b0 : btn_paris_raw; // BTN 5 -> Paris
    wire clk_uk_p    = (sw_alarm) ? 1'b0 : btn_uk_raw;    // BTN 6 -> UK
    
    // �˶� ���� (SW4 ON): ���� ����
    // 4��->�˶�1, 5��->�˶�2, 6��->�˶�3
    wire alm_slot1_p = (sw_alarm) ? btn_ny_raw    : 1'b0; // BTN 4 -> Slot 1
    wire alm_slot2_p = (sw_alarm) ? btn_paris_raw : 1'b0; // BTN 5 -> Slot 2
    wire alm_slot3_p = (sw_alarm) ? btn_uk_raw    : 1'b0; // BTN 6 -> Slot 3


    // ==================================================
    // 2. ���� �ð� ���� 
    // ==================================================
    wire [5:0] wc_sec, wc_min;
    wire [4:0] hour_kst, hour24, hour_disp;
    wire mode_12h, is_pm;
    wire [1:0] tz_sel;

    time_base U_TIME (
        .clk      (clk),
        .rst      (rst),
        .adj_min_p(time_adj_min_p),
        .adj_hour_p(time_adj_hour_p),
        .sec      (wc_sec),
        .min      (wc_min),
        .hour     (hour_kst)
    );

    tz_mode_ctrl U_MODE (
        .clk            (clk),
        .rst            (rst),
        .mode_toggle_p (mode_toggle_p),
        .paris_p        (clk_paris_p), // BTN 5
        .ny_p           (clk_ny_p),    // BTN 4
        .uk_p           (clk_uk_p),    // BTN 6
        .korea_p        (btn_korea_raw),// BTN 7
        .mode_12h       (mode_12h),
        .tz_sel         (tz_sel)
    );

    world_time_calc U_WT (
        .hour_kst(hour_kst),
        .tz_sel  (tz_sel),
        .hour24  (hour24)
    );

    hour12_24 U_HMODE (
        .hour24  (hour24),
        .mode_12h(mode_12h),
        .hour_disp(hour_disp),
        .is_pm   (is_pm)
    );

    wire [3:0] wc_h_ten, wc_h_one;
    wire [3:0] wc_m_ten, wc_m_one;
    wire [3:0] wc_s_ten, wc_s_one;

    hms_to_bcd U_BCD_WC (
        .hour_disp(hour_disp),
        .min      (wc_min),
        .sec      (wc_sec),
        .h_ten    (wc_h_ten), .h_one(wc_h_one),
        .m_ten    (wc_m_ten), .m_one(wc_m_one),
        .s_ten    (wc_s_ten), .s_one(wc_s_one)
    );
    
    // ==================================================
    // [�˶� �ð� ���] - 3 Slot Multi Alarm
    // ==================================================
    wire alarm_ringing;
    wire [3:0] alm_h_ten, alm_h_one;
    wire [3:0] alm_m_ten, alm_m_one;
    wire [2:0] edit_slot; // ���� ���� ���� ���� ��ȣ
    wire a1_en, a2_en, a3_en;
    
    assign alm_led1 = a1_en;
    assign alm_led2 = a2_en;
    assign alm_led3 = a3_en;

    alarm_clock U_ALARM (
        .clk(clk), .rst(rst),
        .sw_alarm(sw_alarm),
        .btn_hour_p(alarm_adj_hour_p),
        .btn_min_p(alarm_adj_min_p),
        .btn_slot1_p(alm_slot1_p), // BTN 4
        .btn_slot2_p(alm_slot2_p), // BTN 5
        .btn_slot3_p(alm_slot3_p), // BTN 6
        .btn_reset_p(btn_alarm_reset_p), // BTN 8 (Reset All - SW3 OFF�϶���)
        .btn_stop_p(alarm_stop_signal),  // *,0,# (Turn Off)
        .curr_hour(hour24),              // 24�ð��� ��
        .curr_min(wc_min),
        .curr_sec(wc_sec),
        .alarm_ringing(alarm_ringing),
        .edit_slot(edit_slot),
        .alm1_en(a1_en), .alm2_en(a2_en), .alm3_en(a3_en),
        .alm_h_ten(alm_h_ten), .alm_h_one(alm_h_one),
        .alm_m_ten(alm_m_ten), .alm_m_one(alm_m_one)
    );

    // ==================================================
    // 3. Ÿ�̸� ���� 
    // ==================================================
    wire [5:0] tm_min_val, tm_sec_val;
    wire tm_alarm;
    wire tm_run_led;
    wire [5:0] tm_init_min_val, tm_init_sec_val; // �ʱ� ���� �ð�

    // [����] Ÿ�̸� ��尡 �����ִ���(SW3 OFF), Ÿ�̸� �˶��� �︮�� ��ư �Է��� ���
    wire tm_min_in   = (sw_timer || tm_alarm) ? tm_min_p : 1'b0;
    wire tm_sec_in   = (sw_timer || tm_alarm) ? tm_sec_p : 1'b0;
    wire tm_start_in = (sw_timer || tm_alarm) ? tm_start_p : 1'b0;

    // [���� 2] Ÿ�̸� ��� �ν��Ͻ� (btn_reset_p �߰� ����)
    timer U_TIMER (
        .clk             (clk),
        .rst             (rst),
        .btn_min_p       (tm_min_in),
        .btn_sec_p       (tm_sec_in),
        .btn_start_stop_p(tm_start_in),
        .btn_reset_p     (btn_timer_reset_p), // SW3 ON�� �� Key 8 �Է�
        .tm_min          (tm_min_val),
        .tm_sec          (tm_sec_val),
        .tm_run_led      (tm_run_led),
        .tm_alarm        (tm_alarm),
        .led_r           (tm_led_r),
        .led_g           (tm_led_g),
        .led_b           (tm_led_b),
        .init_min        (tm_init_min_val),
        .init_sec        (tm_init_sec_val)
    );

    // Ÿ�̸ӿ� BCD ��ȯ
    wire [3:0] tm_m_ten, tm_m_one;
    wire [3:0] tm_s_ten, tm_s_one;

    hms_to_bcd U_BCD_TM (
        .hour_disp(5'd0),
        .min      (tm_min_val),
        .sec      (tm_sec_val),
        .h_ten    (), .h_one(), 
        .m_ten    (tm_m_ten), .m_one(tm_m_one),
        .s_ten    (tm_s_ten), .s_one(tm_s_one)
    );

    // ==================================================
    // 4. ȭ�� ��� ��Ƽ�÷��� (MUX)
    // ==================================================
    wire [3:0] d_h_ten, d_h_one;
    wire [3:0] d_m_ten, d_m_one;
    wire [3:0] d_s_ten, d_s_one;

    // �켱����: SW3(Timer) > SW4(Alarm) > Clock
    assign d_h_ten = sw_timer ? 4'd0 : (sw_alarm ? alm_h_ten : wc_h_ten);
    assign d_h_one = sw_timer ? 4'd0 : (sw_alarm ? alm_h_one : wc_h_one);
    
    assign d_m_ten = sw_timer ? tm_m_ten : (sw_alarm ? alm_m_ten : wc_m_ten);
    assign d_m_one = sw_timer ? tm_m_one : (sw_alarm ? alm_m_one : wc_m_one);
    
    assign d_s_ten = sw_timer ? tm_s_ten : (sw_alarm ? 4'd0 : wc_s_ten); 
    assign d_s_one = sw_timer ? tm_s_one : (sw_alarm ? 4'd0 : wc_s_one);
    
    // DP(�Ҽ���) ����� �߰��� SegDriver
    seg6_driver U_SEG (
        .clk     (clk),
        .rst     (rst),
        .h_ten   (d_h_ten), .h_one(d_h_one),
        .m_ten   (d_m_ten), .m_one(d_m_one),
        .s_ten   (d_s_ten), .s_one(d_s_one),
        .seg_data(seg_data),
        .seg_com (seg_com)
    );

    // ==================================================
    // 5. �ǿ��� ���� (���� Ÿ�� / ��ȭ�� / ������ �и�)
    // ==================================================

    // [���� �˸��� ��������]
    reg hourly_active;      
    reg [3:0] hourly_cnt;   
    reg [3:0] hourly_target;
    reg [9:0] hourly_timer; 
    reg hourly_out;         

    // ��(sec) ��ȭ ���� (���� Ʈ���ſ�)
    reg [5:0] wc_sec_prev;
    always @(posedge clk) wc_sec_prev <= wc_sec;
    wire sec_tick = (wc_sec != wc_sec_prev); // 1�ʿ� �� �� High

    // [��ȭ�� ȿ���� �������� (�˶��ð��)]
    reg [5:0] trill_cnt; 
    reg tone_sel;        
    reg freq_div;        
    
    // [Ÿ�̸ӿ� �߻� ī����]
    reg [9:0] beep_cnt;  

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            piezo <= 0;
            trill_cnt <= 0; tone_sel <= 0; freq_div <= 0;
            beep_cnt <= 0;
            hourly_active <= 0; hourly_cnt <= 0; hourly_target <= 0; hourly_timer <= 0; hourly_out <= 0;
        end else begin
            
            // ----------------------------------------------------
            // A. ���� �˸� ���� (�ð� ����ŭ ��- ��- ��-)
            // ----------------------------------------------------
            if (sec_tick && (wc_min == 0) && (wc_sec == 0)) begin
                hourly_active <= 1;
                hourly_cnt <= 0;
                hourly_timer <= 0;
                hourly_out <= 1; // ��! ����
                
                // Ÿ�� Ƚ�� ��� (12�ð��� ��ȯ)
                if (hour_kst == 0) hourly_target <= 4'd12;               // 0�� -> 12��
                else if (hour_kst <= 12) hourly_target <= hour_kst[3:0]; // 1~12��
                else hourly_target <= hour_kst - 5'd12;                  // 13~23�� -> 1~11��
            end

            if (hourly_active) begin
                if (hourly_timer >= 499) begin
                    hourly_timer <= 0;
                    if (hourly_cnt + 1 >= hourly_target) begin
                        hourly_active <= 0; // ��ǥ Ƚ�� ä��� ����
                        hourly_out <= 0;
                    end else begin
                        hourly_cnt <= hourly_cnt + 1;
                        hourly_out <= 1; // ���� ��! ����
                    end
                end else begin
                    hourly_timer <= hourly_timer + 1;
                    if (hourly_timer < 200) hourly_out <= 1; // 200ms ON
                    else hourly_out <= 0;                    // 300ms OFF
                end
            end else begin
                hourly_out <= 0;
            end

            // ----------------------------------------------------
            // B. ī���� ������Ʈ
            // ----------------------------------------------------
            // �˶��ð�(��ȭ��)�� (50ms �ֱ�)
            if (trill_cnt >= 49) begin
                trill_cnt <= 0; tone_sel <= ~tone_sel;
            end else trill_cnt <= trill_cnt + 1;
            
            freq_div <= ~freq_div; // 250Hz ������ ���� 2����

            // Ÿ�̸ӿ� (0.5�� �ֱ�)
            if (beep_cnt >= 999) beep_cnt <= 0;
            else beep_cnt <= beep_cnt + 1;

            // ----------------------------------------------------
            // C. Piezo ��� MUX (�켱����: �˶��ð� > Ÿ�̸� > ����)
            // ----------------------------------------------------
            if (alarm_ringing) begin
                // [TYPE 1] �˶� �ð�: ��ȭ�� (Trill)
                if (tone_sel == 0) piezo <= ~piezo; // 500Hz
                else if (freq_div) piezo <= ~piezo; // 250Hz
            end
            else if (tm_alarm) begin
                // [TYPE 2] Ÿ�̸�: �ܼ� ��-�� (0.5�� ����)
                if (beep_cnt < 500) piezo <= ~piezo;
                else piezo <= 0;
            end
            else if (hourly_active && hourly_out) begin
                // [TYPE 3] ���� �˸�: ª�� ��! (�ð� ����ŭ �ݺ�)
                piezo <= ~piezo; // 500Hz ��
            end
            else begin
                piezo <= 0;
            end
        end
    end

    // ==================================================
    // 6. LCD ��� �ν��Ͻ� (���� ����)
    // ==================================================
    lcd_worldclock U_LCD (
        .clk(clk), .rst(rst),
        .mode_12h(mode_12h), .tz_sel(tz_sel), .is_pm(is_pm),
        .sw_timer(sw_timer),
        .tm_alarm(tm_alarm),
        .sw_alarm(sw_alarm),
        .alarm_ringing(alarm_ringing),
        
        .edit_slot(edit_slot),
        .alm1_en(a1_en), .alm2_en(a2_en), .alm3_en(a3_en),
        
        .tm_running(tm_run_led), 
        .tm_init_min(tm_init_min_val),
        .tm_init_sec(tm_init_sec_val),
        
        .LCD_E(LCD_E), .LCD_RS(LCD_RS), .LCD_RW(LCD_RW), .LCD_DATA(LCD_DATA)
    );
endmodule